module main

enum TokenKind {
	right_tilde_arrow
	left_tilde_arrow
	plus
	minus
	look
	dollar
	left_brackets
	right_brackets
}
